 
 Timer Timer_inst(
  .CPUdat(CPUdat),
  .CPUctr(CPUctr),

  .Evnt0(Evnt0),
  .Evnt1(Evnt1),
  .Evnt2(Evnt2),
  .PWM(PWM),
	
  .Int(Int),
  .Rst(Rst),
  .Clk(Clk)
 );
